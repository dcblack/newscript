// Project: winnie
// Design:  example
// FILE:   ABOUT_example.txt
/*/////////////////////////////////////////////////////////////////////////
Widgets Inc. PROPRIETARY AND CONFIDENTIAL
Copyright 2010 Widgets Inc..

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

  http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.

/*/////////////////////////////////////////////////////////////////////////
// {:LONG_DESCRIPTION:}
//
// Author :       {:AUTHOR:}
// Contact info : {:EMAIL:}
///////////////////////////////////////////////////////////////////////////
// Version control information
//
// $Source$
// $Id$
// $Revision$
///////////////////////////////////////////////////////////////////////////
//
// {:DUT_DESCRIPTION:}

module widget2_rtl(
( {:DUT_DIR_{:uc:DIR0:}:} {:DUT_TYPE_{:uc:DIR0:}:} [1-1:0] clk
, {:DUT_DIR_{:uc:DIR1:}:} {:DUT_TYPE_{:uc:DIR1:}:} [1-1:0] data_in
, {:DUT_DIR_{:uc:DIR2:}:} {:DUT_TYPE_{:uc:DIR2:}:} [1-1:0] data_out
);

  {:BEHAVIOR_OR_STRUCTURE:}

endmodule
